// MIPS Top Module
// Nicolas Rodriguez
// Nov. 23, 2020

module mips_cpu_revB (clk, reset);

// i/o
input clk, reset;

// local
// assign wires
// combinational logic
// sequential logic
// instances

endmodule // mips_cpu_revB
